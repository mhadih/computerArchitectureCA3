`timescale 1ns/1ns 
module zeroExtend(input [4:0] pc,output [7:0] out);
  assign out = {3'b0,ipc};
endmodule 