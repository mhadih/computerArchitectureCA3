`timescale 1ns/1ns
module DataPath(input clk,rst,
                    pcWrite, pcWriteCond, pcSrc, IorD, memRead, memWrite, IRWrite, MtoS
                    ldA, ldB, srcA, srcB, ALUOp, push, pop, tos
                    input [1:0] func,
                output zero,
                output[2:0] opcode,
                output[4:0] Addrs);
    

endmodule